/*
    This module is used for creating the FIB table of the NDN router. The FIB table consists of 
    
*/

module (
    
);

endmodule // 