module spi_interface_module();

// SPI interfaces
wire sclk;
wire mosi;
reg miso;
wire cs;

// Overall inputs
reg clk;
reg rst;

// Receiving output
wire          RX_valid;  // Valid pulse for 1 cycle for RX byte to know data is ready
wire		  output_shift_register;

// Transferring input
reg               TX_valid;                   // Valid pulse for 1 cycle for TX byte
wire [7:0]        input_shift_register;

reg [1:0] state;
parameter tx = 0, waiting = 1, sending = 2;    

// Instantiate the module
spi_interface spi_interface_module(
    .sclk(sclk),
    .mosi(mosi),
    .miso(miso),
    .cs(cs),
    .clk(clk),
    .rst(rst),
    .RX_valid(RX_valid),
	.output_shift_register(output_shift_register),
    .TX_valid(TX_valid),
	.input_shift_register(input_shift_register)
);

/*
    VALUES USED FOR SIMULATION
*/
reg start_incoming_packet;
reg start_outgoing_packet;

reg [7:0]         packet_meta_data_test;     
reg [71:0]        packet_prefix_test;
reg [255:0]       packet_data_test;
reg [327:0]		  transmitting_data_test;

assign input_shift_register = transmitting_data_test[327:320];

initial begin
    TX_valid = 0;
    start_incoming_packet = 0;
    start_outgoing_packet = 0;
	clk = 0;
    rst = 0;
	state = 0;

    // Start outgoing packet
    packet_meta_data_test = 8'b00101000;
    packet_prefix_test = 64'd129;
    packet_data_test = "here is data";
	transmitting_data_test = {packet_meta_data_test, packet_prefix_test, packet_data_test};
end


always
begin
	// Create clock
	#10 clk = ~clk;
	if(clk) begin
		case(state)
		tx:
		begin
			TX_valid <= 1;
			state <= waiting;
		end
		waiting:
		begin
			TX_valid <= 0;
			state <= sending;
		end
		sending:
		begin
			transmitting_data_test <= transmitting_data_test << 8;
		end
		endcase

	end
end

endmodule
