/*
    This SPI module is used to from NDN --> MCU (user).
    In this set up the NDN module acts as the slave, and the MCU acts as the
    master.
*/
module spi_mcu(
    input sclk,
    input mosi,
    output mosi,
    input ss
);



endmodule 